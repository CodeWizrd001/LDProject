module StimTraffic ;


initial
begin

end
endmodule 