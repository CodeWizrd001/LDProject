module StimTraffic ;

wire [5:0] ans ;
reg clk ;
reg [1023:0] imgData ;
reg [1023:0] Data ;

integer Fin,Fin_ ;

TrafficSystem a(clk,imgData,ans) ;

initial
begin
	clk = 0 ;
end 

always
begin
	clk=~clk ;#1 ;
end

initial
begin
	imgData = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111100000000001111111111111111111111100000000011111111111111111111111000000000000000000000000001111100000000000000000000000000011111000000000000000000000000000111110000000000000000000000000111111000000000000000000000000001111100000000000000000000000000111110000000000000000000000000111111000000000000000000000000001111100000000000000000000000000111111000000000000000000000000011111000000000000000000000000000111110000000000000000000000000111111000000000000000000000000001111110000000000000000000000000111110000000000000000000000000001111100000000000000000000000000111110000000000000000000000000111111000000000000000000000000001111110000000000000000000000000111110000000000000000000000000001111000000000000000000000000000111110000000000000000000000000111111000000000000000000000000001111000000000000000000000000000011110000000000000000000000000001111111111111111111111110000000011111111111111111111111100000000011111111111111111111111000 ; #5 ;
	imgData = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000001111111111111000000000000000000011111111111111000000000000000000111000000011111000000000000000001110000000011110000000000000000011100000000011110000000000000000111000000000111100000000000000001110000000001111000000000000000011100000000011110000000000000000111000000000111000000000000000001110000000011110000000000000000011100000001111000000000000000000111111111111100000000000000000001111111111111000000000000000000011111111111111100000000000000000111000000001111100000000000000001110000000000111100000000000000011100000000001111000000000000000111000000000001110000000000000001110000000000011100000000000000011100000000000111000000000000000111000000000011110000000000000001110000000000111100000000000000011100000000111110000000000000000111111111111111000000000000000001111111111111100000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ; #5 ; 
	imgData = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000111111111110000000000000000000011111111111111000000000000000001111100000011110000000000000000111100000000001110000000000000011110000000000001100000000000000111100000000000000000000000000011110000000000000000000000000000111100000000000000000000000000001110000000000000000000000000000111100000000000000000000000000001111000000000000000000000000000011110000000000000000000000000000111100000000000000000000000000001111000000000000000000000000000011110000000000000000000000000000111100000000000000000000000000001111000000000000000000000000000001111000000000000000000000000000011110000000000000000000000000000111100000000000000000000000000000111100000000000011000000000000001111100000000001110000000000000001111110000001111100000000000000001111111111111110000000000000000000111111111110000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ; #5 ;
	$system("python ProcessImage.py A_1") ; #5 ;
	Fin = $fopen("A_0.txt","r") ;
	Fin_ = $fscanf(Fin,"%b",imgData) ; #5 ;
end
endmodule 